module immSrcControl(input [1:0] opType,output immSrc);

	assign immSrc= opType[0];
endmodule 